


 package router_test_pkg;




import uvm_pkg::*;


`include "uvm_macros.svh"


`include "typedefs.sv"

`include "src_xtns.sv"
`include "src_agent_config.sv"
`include "dst_agent_config.sv"
`include "src_seq.sv"
`include "env_config.sv"
`include "src_driver.sv"
`include "src_sequencer.sv"
`include "src_monitor.sv"
`include "src_agent.sv"
`include "src_top.sv"



`include "dst_xtns.sv"
`include "dst_sequencer.sv"
`include "dst_seqs.sv"
`include "dst_driver.sv"
`include "dst_monitor.sv"
`include "dst_agent.sv"
`include "dst_top.sv"

`include "virtual_sequencer.sv"
`include "virtual_seq.sv"

`include "scoreboard.sv"

`include "router_tb.sv"

`include "test_top.sv"











endpackage
