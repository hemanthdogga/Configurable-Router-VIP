



typedef enum {GOOD_PARITY,BAD_PARITY} parity_type;
